library verilog;
use verilog.vl_types.all;
entity Tb_Adder0 is
end Tb_Adder0;
