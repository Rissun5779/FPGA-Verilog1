module Adder0(
  input  bit x,
  input  bit y,
  input  bit Cin,
  
  output bit Cout,
  output bit Sum
);
  assign {Cout, Sum} = x+y+Cin;
endmodule 